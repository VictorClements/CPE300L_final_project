module numberInputFSM(input  logic clk, reset,
                      input  logic 
);
  
endmodule